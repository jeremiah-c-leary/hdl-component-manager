This would be the rook entity.
