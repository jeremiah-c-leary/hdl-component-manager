This would be a VHDL entity.
