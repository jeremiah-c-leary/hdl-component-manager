This is an extra file that is not in the manifest.
